`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 11/16/2017 02:42:40 PM
// Design Name: 
// Module Name: TopLevel_tb_custom_testcases_1
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module TopLevel_tb_custom_testcases_1();
    
    reg Clk, Rst;
        
    wire [31:0] WriteData, PCValue, HiReg, LoReg;
    
    integer tests, passed;
    
    TopLevel m0(
        .Clk(Clk),
        .Rst(Rst),
        .WriteData(WriteData),
        .PCValue(PCValue),
        .HiReg(HiReg),
        .LoReg(LoReg)
    );
          
    initial begin
        Clk <= 1'b0;
        forever #100 Clk <= ~Clk;
    end
    
    initial begin
        tests <= 0;
        passed <= 0;
        Rst <= 1;
        
        $display("\n\n~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~");
        $display("Starting Unit Tests.");
        
        @(negedge Clk);
        @(negedge Clk);
        Rst <= 0;
        @(negedge Clk);
        @(negedge Clk);
        @(negedge Clk);
        
        // main:
        
        
        // la $s1, asize0        
        @(negedge Clk);
        tests = tests + 1; // Test #1
        #5 if (WriteData == 32'h0)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #1: la $s1, asize0. Exceptect WriteData: 0. Actual WriteData: %h", $time, WriteData);
        
        
        //// BEGIN FORWARDING TESTS ////
        
        
        //// forward to lw address ////
        
        // la $t1, asize0          
        @(negedge Clk);
        tests = tests + 1; // Test #2
        #5 if (WriteData == 32'h0)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #2: la $t1, asize0. Exceptect WriteData: 0. Actual WriteData: %h", $time, WriteData);
        
        // addi $t2, $t1, 0        
        @(negedge Clk);
        tests = tests + 1; // Test #3
        #5 if (WriteData == 32'h0)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #3: addi $t2, $t1, 0. Exceptect WriteData: 0. Actual WriteData: %h", $time, WriteData);
        
        // lw $t3, 4($t2)          
        @(negedge Clk);
        tests = tests + 1; // Test #4
        #5 if (WriteData == 32'd200)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #4: lw $t3, 4($t2). Exceptect WriteData: 200. Actual WriteData: %d", $time, WriteData);
        
        
        //// forward to sw address ////
        
        // addi $t4, $zero, 5      
        @(negedge Clk);
        tests = tests + 1; // Test #5
        #5 if (WriteData == 32'd5)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #5: addi $t4, $zero, 5. Exceptect WriteData: 5. Actual WriteData: %d", $time, WriteData);
        
        // add $t3, $zero, $t1     
        @(negedge Clk);
        tests = tests + 1; // Test #6
        #5 if (WriteData == 32'h0)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #6: add $t3, $zero, $t1. Exceptect WriteData: 0. Actual WriteData: %h", $time, WriteData);
        
        // sw $t4, 4($t3)
        @(negedge Clk);
        
        // lw $t2, 4($t3)          
        @(negedge Clk);
        tests = tests + 1; // Test #7
        #5 if (WriteData == 32'd5)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #7: lw $t2, 4($t3). Exceptect WriteData: 5. Actual WriteData: %d", $time, WriteData);
        
        
        //// sw after lw rt dependency ////
        
        // lw $t1, 0($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #8
        #5 if (WriteData == 32'd100)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #8: lw $t1, 0($s1). Exceptect WriteData: 100. Actual WriteData: %d", $time, WriteData);
        
        // sw $t1, 4($s1)
        @(negedge Clk);
        
        // lw $t2, 4($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #9
        #5 if (WriteData == 32'd100)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #9: lw $t2, 4($s1). Exceptect WriteData: 100. Actual WriteData: %d", $time, WriteData);
        
        
        //// sw after add rt dependency ////
        
        // add $t1, $t1, $t1       
        @(negedge Clk);
        tests = tests + 1; // Test #10
        #5 if (WriteData == 32'd200)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #10: add $t1, $t1, $t1. Exceptect WriteData: 200. Actual WriteData: %d", $time, WriteData);
        
        // sw $t1, 8($s1)
        @(negedge Clk);
        
        // lw $t3, 8($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #11
        #5 if (WriteData == 32'd200)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #11: lw $t3, 8($s1). Exceptect WriteData: 200. Actual WriteData: %d", $time, WriteData);
        
        
        //// sw after unrelated after lw dependency ////
        
        // lw $t3, 12($s1)         
        @(negedge Clk);
        tests = tests + 1; // Test #12
        #5 if (WriteData == 32'd400)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #12: lw $t3, 12($s1). Exceptect WriteData: 400. Actual WriteData: %d", $time, WriteData);
        
        // addi $s2, $zero, 15     
        @(negedge Clk);
        tests = tests + 1; // Test #13
        #5 if (WriteData == 32'd15)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #13: addi $s2, $zero, 15. Exceptect WriteData: 15. Actual WriteData: %d", $time, WriteData);
        
        // sw $t3, 16($s1)
        @(negedge Clk);
        
        // lw $t4, 16($s1)         
        @(negedge Clk);
        tests = tests + 1; // Test #14
        #5 if (WriteData == 32'd400)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #14: lw $t4, 16($s1). Exceptect WriteData: 400. Actual WriteData: %d", $time, WriteData);
        
        
        //// sw after unrelated after add dependency ////
        
        // addi $t5, $zero, 7      
        @(negedge Clk);
        tests = tests + 1; // Test #15
        #5 if (WriteData == 32'd7)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #15: addi $t5, $zero, 7. Exceptect WriteData: 7. Actual WriteData: %d", $time, WriteData);
        
        // add $t6, $t5, $t5       
        @(negedge Clk);
        tests = tests + 1; // Test #16
        #5 if (WriteData == 32'd14)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #16: add $t6, $t5, $t5. Exceptect WriteData: 14. Actual WriteData: %d", $time, WriteData);
        
        // sw $t5, 0($s1)
        @(negedge Clk);
        
        // lw $t6, 0($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #17
        #5 if (WriteData == 32'd7)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #17: lw $t6, 0($s1). Exceptect WriteData: 7. Actual WriteData: %d", $time, WriteData);
        
        
        //// r-type after mfhi ////
        
        // mthi $t5
        @(negedge Clk);
        
        // mfhi $t7                
        @(negedge Clk);
        tests = tests + 1; // Test #18
        #5 if (WriteData == 32'd7)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #18: mfhi $t7. Exceptect WriteData: 7. Actual WriteData: %d", $time, WriteData);
        
        // ori $s2, $t7, 8         
        @(negedge Clk);
        tests = tests + 1; // Test #19
        #5 if (WriteData == 32'd15)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #19: ori $s2, $t7, 8. Exceptect WriteData: 15. Actual WriteData: %d", $time, WriteData);
        
        
        //// r-type after mflo ////
        
        // mtlo $t3
        @(negedge Clk);
        
        // mflo $s2                
        @(negedge Clk);
        tests = tests + 1; // Test #20
        #5 if (WriteData == 32'd400)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #20: mflo $s2. Exceptect WriteData: 400. Actual WriteData: %d", $time, WriteData);
        
        // slt $s3, $t6, $s2       
        @(negedge Clk);
        tests = tests + 1; // Test #21
        #5 if (WriteData == 32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #21: slt $s3, $t6, $s2. Exceptect WriteData: 1. Actual WriteData: %d", $time, WriteData);
        
        
        //// sw after unrelated after mflo ////
        
        // mflo $s3                
        @(negedge Clk);
        tests = tests + 1; // Test #22
        #5 if (WriteData == 32'd400)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #22: mflo $s3. Exceptect WriteData: 400. Actual WriteData: %d", $time, WriteData);
        
        // addi $s4, $zero, 4      
        @(negedge Clk);
        tests = tests + 1; // Test #23
        #5 if (WriteData == 32'd4)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #23: addi $s4, $zero, 4. Exceptect WriteData: 4. Actual WriteData: %d", $time, WriteData);
        
        // sw $s3, 0($s1)
        @(negedge Clk);
        
        // lw $s4, 0($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #24
        #5 if (WriteData == 32'd400)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #24: lw $s4, 0($s1). Exceptect WriteData: 400. Actual WriteData: %d", $time, WriteData);
        
        
        //// branch after unrelated after r-type ////
        
        // addi $s2, $zero, -1     
        @(negedge Clk);
        tests = tests + 1; // Test #25
        #5 if (WriteData == -32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #25: addi $s2, $zero, -1. Exceptect WriteData: -1. Actual WriteData: %d", $time, WriteData);
        
        // addi $s4, $zero, 4      
        @(negedge Clk);
        tests = tests + 1; // Test #26
        #5 if (WriteData == 32'd4)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #26: addi $s4, $zero, 4. Exceptect WriteData: 4. Actual WriteData: %d", $time, WriteData);
        
        // bgez $s2, error         
        @(negedge Clk);
        
        // addi $s5, $zero, 5      
        @(negedge Clk);
        tests = tests + 1; // Test #27
        #5 if (WriteData == 32'd5)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #27: addi $s5, $zero, 5. Exceptect WriteData: 5. Actual WriteData: %d", $time, WriteData);
        
        
        //// branch after unrelated after r-type 2 ////
        
        // add $s6, $zero, $s5    
        @(negedge Clk);
        tests = tests + 1; // Test #28
        #5 if (WriteData == 32'd5)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #28: addi $s6, $zero, $s5. Exceptect WriteData: 5. Actual WriteData: %d", $time, WriteData);
        
        // addi $s4, $zero, 3      
        @(negedge Clk);
        tests = tests + 1; // Test #29
        #5 if (WriteData == 32'd3)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #29: addi $s4, $zero, 3. Exceptect WriteData: 3. Actual WriteData: %d", $time, WriteData);
        
        // beq $s5, $s6, branch1   
        @(negedge Clk);
        
        // Flush 
        @(negedge Clk);
        
        // branch1:
        
        // addi $s5, $zero, 1      
        @(negedge Clk);
        tests = tests + 1; // Test #30
        #5 if (WriteData == 32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #30: addi $s5, $zero, 1. Exceptect WriteData: 1. Actual WriteData: %d", $time, WriteData);
        
        
        //// branch after unrelated after mfhi ////
        
        // mfhi $s4                
        @(negedge Clk);
        tests = tests + 1; // Test #31
        #5 if (WriteData == 32'd7)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #31: mfhi $s4. Exceptect WriteData: 7. Actual WriteData: %d", $time, WriteData);
        
        // addi $s5, $zero, 2      
        @(negedge Clk);
        tests = tests + 1; // Test #32
        #5 if (WriteData == 32'd2)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #32: addi $s5, $zero, 2. Exceptect WriteData: 2. Actual WriteData: %d", $time, WriteData);
        
        // bgtz $s4, branch2       
        @(negedge Clk);
        
        // Flush
        @(negedge Clk);
        
        // branch2:
        
        // addi $s5, $zero, 1      
        @(negedge Clk);
        tests = tests + 1; // Test #33
        #5 if (WriteData == 32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #33: addi $s5, $zero, 1. Exceptect WriteData: 1. Actual WriteData: %d", $time, WriteData);
        
        
        //// BEGIN STALLING TESTS ////
        
        // la $s1, asize1
        @(negedge Clk);
        
        // sw $s1, 0($s1)
        @(negedge Clk);
        
        
        //// sw after lw ////
        
        // lw $s2, 0($s1)
        @(negedge Clk);
        
        // Stalling. 
        @(negedge Clk);
        
        // sw $s5, 4($s2)
        @(negedge Clk);
        
        // lw $s6, 4($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #34
        #5 if (WriteData == 32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #34: lw $s6, 4($s1). Exceptect WriteData: 1. Actual WriteData: %d", $time, WriteData);
        
        
        //// r-type after lw ////
        
        // Stalling. 
        @(negedge Clk);
        
        // add $s5, $s6, $s6       
        @(negedge Clk);
        tests = tests + 1; // Test #35
        #5 if (WriteData == 32'd2)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #35: add $s5, $s6, $s6. Exceptect WriteData: 2. Actual WriteData: %d", $time, WriteData);
        
        
        //// branch after r-type ////
        
        // addi $s5, $zero, -3     
        @(negedge Clk);
        tests = tests + 1; // Test #36
        #5 if (WriteData == -32'd3)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #36: addi $s5, $zero, -3. Exceptect WriteData: -3. Actual WriteData: %d", $time, WriteData);
        
        // Stalling. 
        @(negedge Clk);
        
        // bgez $s5, error         
        @(negedge Clk);
        
        // addi $s2, $zero, -1      
        @(negedge Clk);
        tests = tests + 1; // Test #37
        #5 if (WriteData == -32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #37: addi $s2, $zero, -1. Exceptect WriteData: -1. Actual WriteData: %d", $time, WriteData);
        
        
        //// branch after lw ////
        
        // lw $s2, 8($s1)          
        @(negedge Clk);
        tests = tests + 1; // Test #38
        #5 if (WriteData == 32'd900)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #38: lw $s2, 8($s1). Exceptect WriteData: 900. Actual WriteData: %d", $time, WriteData);
        
        // Stalling. 
        @(negedge Clk);
        
        // Stalling. 
        @(negedge Clk);
        
        // bgez $s2, branch3       
        @(negedge Clk);
        
        // Flush
        @(negedge Clk);
        
        // branch3:
        
        // addi $s2, $zero, 1      
        @(negedge Clk);
        tests = tests + 1; // Test #39
        #5 if (WriteData == 32'd1)
            passed = passed + 1;
        else
            $display("Time: %0d. Failed Test #39: addi $s2, $zero, 1. Exceptect WriteData: 1. Actual WriteData: %d", $time, WriteData);
        
        // done:
        
        // j done
        @(negedge Clk);
        
        // Report results
        if (passed == tests)
            $display("All tests passed.");
        else
            $display("%3d out of %3d tests passed.", passed, tests);
        $display("~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~~\n\n");

    end
endmodule
