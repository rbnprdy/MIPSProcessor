`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// ECE369A - Computer Architecture
// Laboratory  1
// Module - InstructionMemory.v
// Description - 32-Bit wide instruction memory.
//
// INPUT:-
// Address: 32-Bit address input port.
//
// OUTPUT:-
// Instruction: 32-Bit output port.
//
// FUNCTIONALITY:-
// Similar to the DataMemory, this module should also be byte-addressed
// (i.e., ignore bits 0 and 1 of 'Address'). All of the instructions will be 
// hard-coded into the instruction memory, so there is no need to write to the 
// InstructionMemory.  The contents of the InstructionMemory is the machine 
// language program to be run on your MIPS processor.
//
//
//we will store the machine code for a code written in C later. for now initialize 
//each entry to be its index * 4 (memory[i] = i * 4;)
//all you need to do is give an address as input and read the contents of the 
//address on your output port. 
// 
//Using a 32bit address you will index into the memory, output the contents of that specific 
//address. for data memory we are using 1K word of storage space. for the instruction memory 
//you may assume smaller size for practical purpose. you can use 128 words as the size and 
//hardcode the values.  in this case you need 7 bits to index into the memory. 
//
//be careful with the least two significant bits of the 32bit address. those help us index 
//into one of the 4 bytes in a word. therefore you will need to use bit [8-2] of the input address. 


////////////////////////////////////////////////////////////////////////////////

module InstructionMemory(Address, Instruction); 

    input [31:0] Address;        // Input Address 

    output reg [31:0] Instruction;    // Instruction at memory location Address
    
    reg [31:0] memory [0:395]; // memory is an array with 9 32 bit numbers ([lsb:msb] is convention for words)
    
    initial begin
        //$readmemh("C:/Users/Ruben Purdy/Documents/ECE369/processor/Instruction_memory_custom_testcases_jump.txt", memory); // place "Instruction_memory.txt" in PROJECT_NAME.sim\sim_1\behav\xsim  
        memory[0] = 32'b00100000000010000000000000000101; // addi $t0, $zero, 5
        memory[1] = 32'b00001100000000000000000000000101; // jal 5
        memory[2] = 32'b00100000000010000000000000000101; // addi $t0, $zero, 6
        memory[3] = 32'b00100000000010000000000000000111; // addi $t0, $zero, 7
        memory[4] = 32'b00100000000010000000000000001000; // addi $t0, $zero, 8
        memory[5] = 32'b00100000000010000000000000001001; // addi $t0, $zero, 9
        memory[6] = 32'b00100000000010000000000000001010; // addi $t0, $zero, 10
        memory[7] = 32'b00000011111000000000000000001000; // jr $ra
        memory[8] = 32'b00100000000010000000000000001011; // addi $t0, $zero, 11
    end
    
    always @(Address) begin
        Instruction <= memory[Address[10:2]]; // Assign the instruction at the byte address of Address.
    end   

endmodule
